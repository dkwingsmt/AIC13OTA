.param input_diff=1.127831