.param input_diff=0.663796