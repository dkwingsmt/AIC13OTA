.param ib=2.0691e-04
.param cl=3.9962e-12
.param cs=4.0000e-12
.param cf=2.0000e-12
.param ln=4.1017e-07
.param lp=6.3338e-07
.param wb=2.1964e-05
.param w0=4.3928e-04
.param w1=8.1734e-04
.param w2=8.1734e-04
.param w1a=2.1623e-04
.param w2a=2.1623e-04
.param w3=1.1957e-03
.param w3a=1.1957e-03
.param w4=1.1957e-03
.param w4a=1.1957e-03
.param w5a=5.0221e-05
.param w5b=2.5110e-04
.param w5c=4.3928e-05
.param w6a=1.1957e-04
.param w6b=1.1957e-04
.param w6c=1.7298e-05
.param w6d=3.4597e-06
.param w7a=2.5110e-04
.param w7b=2.5110e-04
.param w7c=4.3928e-05
