.param input_diff=0.824603