.param input_diff=0.822167