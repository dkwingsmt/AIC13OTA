.param ib=2.0691e-04
.param cl=2.3000e-12
.param cs=6.6000e-12
.param cf=3.3000e-12
.param ln=4.1017e-07
.param lp=6.3338e-07
.param wb=2.1964e-05
.param w0=4.3928e-04
.param w1=6.5387e-04
.param w2=6.5387e-04
.param w1a=3.2434e-04
.param w2a=3.2434e-04
.param w3=1.6142e-03
.param w3a=8.3701e-04
.param w4=1.6142e-03
.param w4a=8.3701e-04
.param w5a=1.7577e-05
.param w5b=8.7886e-05
.param w5c=2.1964e-05
.param w6a=1.6142e-04
.param w6b=8.3701e-05
.param w6c=3.2434e-05
.param w6d=6.4868e-06
.param w7a=1.6949e-04
.param w7b=1.6949e-04
.param w7c=2.1964e-05
.param l12=4.1017e-07
.param l1a=5.3322e-07
.param l3a=6.3338e-07
.param l3=8.5506e-07
.param lbb1p=6.3338e-07
.param lbiasp=6.3338e-07
.param lbb2p1=6.3338e-07
.param lbb2p2=6.3338e-07
.param lbb2n=5.3322e-07
