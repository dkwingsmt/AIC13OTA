.param input_diff=0.784862