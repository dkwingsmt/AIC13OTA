.param ib=9.0075e-05
.param cl=3.9962e-12
.param cs=4.0000e-12
.param cf=2.0000e-12
.param ln=4.1017e-07
.param lp=6.3338e-07
.param wb=9.5616e-06
.param w0=1.9123e-04
.param w1=1.0928e-03
.param w2=1.0928e-03
.param w1a=6.8059e-04
.param w2a=6.8059e-04
.param w3=4.9688e-04
.param w3a=4.9688e-04
.param w4=4.9688e-04
.param w4a=4.9688e-04
.param w5a=1.0931e-04
.param w5b=5.4656e-04
.param w5c=9.5616e-05
.param w6a=9.9375e-05
.param w6b=9.9375e-05
.param w6c=1.0889e-04
.param w6d=2.1779e-05
.param w7a=5.4656e-04
.param w7b=5.4656e-04
.param w7c=9.5616e-05
