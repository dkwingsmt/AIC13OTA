.param input_diff=0.791287