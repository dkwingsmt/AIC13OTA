.param input_diff=0.572422