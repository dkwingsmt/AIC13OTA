.param input_diff=0.684155