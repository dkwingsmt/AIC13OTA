.param ib=2.0691e-04
.param cl=2.0000e-12
.param cs=6.0000e-12
.param cf=3.0000e-12
.param ln=4.1017e-07
.param lp=6.3338e-07
.param wb=2.1964e-05
.param w0=4.3928e-04
.param w1=6.5387e-04
.param w2=6.5387e-04
.param w1a=2.8110e-04
.param w2a=2.8110e-04
.param w3=1.6381e-03
.param w3a=1.1957e-03
.param w4=1.6381e-03
.param w4a=1.1957e-03
.param w5a=2.5110e-05
.param w5b=1.2555e-04
.param w5c=2.1964e-05
.param w6a=1.6381e-04
.param w6b=1.1957e-04
.param w6c=2.8110e-05
.param w6d=5.6219e-06
.param w7a=1.7201e-04
.param w7b=1.7201e-04
.param w7c=2.1964e-05
.param l12=4.5119e-07
.param l1a=4.9220e-07
.param l3a=6.3338e-07
.param l3=8.6773e-07
.param lbb1p=6.3338e-07
.param lbiasp=6.3338e-07
.param lbb2p1=6.3338e-07
.param lbb2p2=6.3338e-07
.param lbb2n=4.9220e-07
