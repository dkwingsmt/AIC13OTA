.param l3=4.0000e-07
.param ib=1.2277e-04
.param cl=5.0955e-12
.param cs=4.0000e-12
.param cf=2.0000e-12
.param ln=4.2670e-07
.param lp=6.2672e-07
.param wb=4.7832e-05
.param w0=9.5663e-04
.param w1=1.1485e-03
.param w2=1.1485e-03
.param w1a=1.0475e-03
.param w2a=1.0475e-03
.param w3=8.3726e-04
.param w3a=8.3726e-04
.param w4=8.3726e-04
.param w4a=8.3726e-04
.param w5a=2.0094e-04
.param w5b=1.0047e-03
.param w5c=4.7832e-04
.param w6a=3.3490e-04
.param w6b=3.3490e-04
.param w6c=3.3519e-04
.param w6d=6.7038e-05
.param w7a=1.0047e-03
.param w7b=1.0047e-03
.param w7c=4.7832e-04
