.param input_diff=0.542309