.param input_diff=0.805265