.param input_diff=0.613742