.param input_diff=0.648216