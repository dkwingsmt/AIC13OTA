.param ib=2.4700e-04
.param cl=5.0955e-12
.param cs=4.0000e-12
.param cf=2.0000e-12
.param ln=4.3244e-07
.param lp=6.3774e-07
.param wb=2.6219e-05
.param w0=5.2438e-04
.param w1=8.1302e-04
.param w2=8.1302e-04
.param w1a=7.6840e-04
.param w2a=7.6840e-04
.param w3=1.3625e-03
.param w3a=1.3625e-03
.param w4=1.3625e-03
.param w4a=1.3625e-03
.param w5a=2.9975e-04
.param w5b=1.4987e-03
.param w5c=2.6219e-04
.param w6a=2.7250e-04
.param w6b=2.7250e-04
.param w6c=1.2294e-04
.param w6d=2.4589e-05
.param w7a=1.4987e-03
.param w7b=1.4987e-03
.param w7c=2.6219e-04
