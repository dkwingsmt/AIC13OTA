.param ib=2.0691e-04
.param cl=3.9962e-12
.param cs=4.0000e-12
.param cf=2.0000e-12
.param ln=4.1017e-07
.param lp=6.3338e-07
.param wb=2.1964e-05
.param w0=4.3928e-04
.param w1=8.1734e-04
.param w2=8.1734e-04
.param w1a=4.3246e-04
.param w2a=4.3246e-04
.param w3=1.1957e-03
.param w3a=1.1957e-03
.param w4=1.1957e-03
.param w4a=1.1957e-03
.param w5a=2.5110e-05
.param w5b=1.2555e-04
.param w5c=2.1964e-05
.param w6a=1.1957e-04
.param w6b=1.1957e-04
.param w6c=4.3246e-05
.param w6d=8.6491e-06
.param w7a=1.2555e-04
.param w7b=1.2555e-04
.param w7c=2.1964e-05
.param l12=4.1017e-07
.param l1a=6.5627e-07
.param l3a=8.8673e-07
.param l3=6.3338e-07
.param lbb1p=8.8673e-07
.param lbiasp=7.6006e-07
.param lbb2p1=7.6006e-07
.param lbb2p2=8.8673e-07
.param lbb2n=6.5627e-07
